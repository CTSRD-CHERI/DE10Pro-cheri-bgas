import IOCapAxi_KeyManager2s :: *;
import IOCapAxi_Exposers_V6 :: *;
import IOCapAxi_Checker3s :: *;
import BlueBasics :: *;
import Tests :: *;
import IOCapAxi_Konata :: *;

// HACK: implement a zero-sized pool (to see the fmax and size for only the surrounding HW) by implementing the Checkers as null variants
(* synthesize *)
module mkCombinedIOCapExposerV6_0pool_1percycle_KeyManager2V1_Tb(UnifiedSingleExposerKeyMngrTb);
    NumProxy#(1) exposerPoolSize = ?;

    let keyMgr32Impl <- mkIOCapAxi_KeyManager2_V1;
    let exposerImpl <- mkSimpleIOCapExposerV6(
        KONATA_FLIT, keyMgr32Impl.exposerPorts[0], True,
        exposerPoolSize,
        mkNullIOCapAxiChecker3V1_Read,
        mkNullIOCapAxiChecker3V1_Write
    );

    interface keyStore = keyMgr32Impl.hostFacingSlave;
    interface debugKeyState = keyMgr32Impl.debugKeyState;
    interface debugGoodWrite = keyMgr32Impl.debugGoodWrite;
    interface debugBadWrite = keyMgr32Impl.debugBadWrite;
    interface debugGoodRead = keyMgr32Impl.debugGoodRead;
    interface debugBadRead = keyMgr32Impl.debugBadRead;
    interface exposer4x32 = exposerImpl;
endmodule